module distancias();

endmodule