//unidade responsável por traduzir os dados para enviar e receber do esp