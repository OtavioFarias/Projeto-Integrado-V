module mapas #(parameter int TamanhoMalha = 20, parameter int tamanhoDistancia = 8 /* em bits*/)(

	input clock,
	input reset,
	
	input [tamanhoDistancia] posicaoAtualnoEixoX,
	input [tamanhoDistancia] posicaoAtualnoEixoY,
	input direcaoAtual, // 0 - horizontal, 1 - vertical
	
	input [tamanhoDistancia] distanciaFrente,
	input [tamanhoDistancia] distanciaDireita,
	input [tamanhoDistancia] distanciaEsquerda,
	
	input novoDado,
	
	
	output reg [1:0] malha[TamanhoMalha][TamanhoMalha], //x,y - 00 - desconhecido, 01 - livre, 10 - ocupado
	output reg operacaoFinalizada // valor 1 se operação finalizada e disponível para receber novas requisições

);

int x,y;

localparam marcarVertical = 2'b00,
		   marcarHorizontal = 2'b01,
		   IDLE = 2'b10;

reg [tamanhoDistancia] marcarDireita;
reg [tamanhoDistancia] marcarEsquerda;

reg [tamanhoDistancia] posicaoDireita;
reg [tamanhoDistancia] posicaoEsquerda;

reg direitaAcabou;
reg esquerdaAcabou;

reg [1:0] stage;

wire [tamanhoDistancia] posicaoEsquerdaX;
wire [tamanhoDistancia] posicaoEsquerdaY;

wire [tamanhoDistancia] posicaoDireitaX;
wire [tamanhoDistancia] posicaoDireitaY;

assign posicaoEsquerdaX = posicaoAtualnoEixoX - distanciaEsquerda;
assign posicaoEsquerdaY = posicaoAtualnoEixoY - distanciaEsquerda;
assign posicaoDireitaX = posicaoAtualnoEixoX + distanciaDireita;
assign posicaoDireitaY = posicaoAtualnoEixoY + distanciaDireita;


always_ff @(posedge clock, posedge reset) begin

	if(reset) begin
	
		 for (x = 0; x < TamanhoMalha; x++) begin
		 	for (y = 0; y < TamanhoMalha; y++) begin
		 
		 		malha[x][y] <= 2'b00;
		 	
		 	end
		 end
		 
		 operacaoFinalizada <= 1'b1;
		 stage <= IDLE;
		 
		marcarDireita <= 0;
		marcarEsquerda <= 0;
		
		direitaAcabou <= 1'b0;
		esquerdaAcabou <= 1'b0;
		 
		posicaoDireita <= 0;
		posicaoEsquerda <= 0;
		 
	end
	else begin
		
		case(stage) 
	
		IDLE: begin
			
			if(novoDado) begin
			
				operacaoFinalizada <= 1'b0;
				
				//marca posição atual
				malha[posicaoAtualnoEixoX][posicaoAtualnoEixoY] <= 2'b01;
				
				// mandar dados para a unidade responsável por marcar
				// aqui os conceitos de direita e esquerda são em relação a posição atual do carrinho
				if(direcaoAtual) begin // vertical be

					marcarDireita  <=  posicaoDireitaX - 1;
					marcarEsquerda <= posicaoEsquerdaX + 1;
					
					// posições atuais da célula a ser marcada, começa na posição atual do carrinho e direciona para até a célula destino
					posicaoDireita <= posicaoAtualnoEixoX;
					posicaoEsquerda <= posicaoAtualnoEixoX;
					
					stage <= marcarVertical;
					
					malha[posicaoDireitaX][posicaoAtualnoEixoY] <= 2'b10;
					malha[posicaoEsquerdaX][posicaoAtualnoEixoY] <= 2'b10;
				
				end
				else begin
				
					marcarDireita  <= posicaoDireitaY - 1;
					marcarEsquerda <= posicaoEsquerdaY + 1;
				
					stage <= marcarHorizontal;
					
					malha[posicaoAtualnoEixoX][posicaoDireitaY] <= 2'b10;
					malha[posicaoAtualnoEixoX][posicaoEsquerdaY] <= 2'b10;
				
					// posições atuais da célula a ser marcada, começa na célula destino e vai até a posição atual do carrinho
					posicaoDireita <= posicaoAtualnoEixoX + distanciaDireita;
					posicaoEsquerda <= posicaoAtualnoEixoX - distanciaEsquerda;
				
				end
			end
			else begin
			
				stage <= IDLE;
			
			end
		end

		marcarHorizontal: begin

			if(direitaAcabou && esquerdaAcabou) begin
			
				direitaAcabou <= 1'b0;
				esquerdaAcabou <= 1'b0;
				
				operacaoFinalizada <= 1'b1;
				
				stage <= IDLE;
			
			end
			else begin 
			
				stage <= marcarHorizontal;

				if(posicaoDireita != marcarDireita) begin

					posicaoDireita  <= posicaoDireita + 1;
					
					malha[posicaoDireita][posicaoAtualnoEixoY] <= 2'b01;
					
				end
				else begin
				
					direitaAcabou <= 1'b1;
				
				end
				
				if(posicaoEsquerda != marcarEsquerda) begin
				
					posicaoEsquerda <= posicaoEsquerda - 1;
					
					malha[posicaoEsquerda][posicaoAtualnoEixoX] <= 2'b01;
				
				end
				else begin
				
					esquerdaAcabou <= 1'b1;
				
				end
			
			end
		end			

		
		marcarVertical: begin
		
			if(direitaAcabou && esquerdaAcabou) begin
			
				direitaAcabou <= 1'b0;
				esquerdaAcabou <= 1'b0;
				
				operacaoFinalizada <= 1'b1;
				
				stage <= IDLE;
			
			end
			else begin 
			
				stage <= marcarVertical;

				if(posicaoDireita != marcarDireita) begin

					posicaoDireita  <= posicaoDireita + 1;
					
					malha[posicaoDireita][posicaoAtualnoEixoY] <= 2'b01;
					
				end
				else begin
				
					direitaAcabou <= 1'b1;
				
				end
				
				if(posicaoEsquerda != marcarEsquerda) begin
				
					posicaoEsquerda <= posicaoEsquerda - 1;
					
					malha[posicaoEsquerda][posicaoAtualnoEixoY] <= 2'b01;
				
				end
				else begin
				
					esquerdaAcabou <= 1'b1;
				
				end
			
			end
		
		end
		
	endcase

				
	end
end

endmodule